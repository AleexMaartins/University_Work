library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

entity TriangSignal_ROM_256x8 is
   port(address : in  std_logic_vector(7 downto 0);
        dataOut : out std_logic_vector(7 downto 0));
end TriangSignal_ROM_256x8;

architecture Behavioral of TriangSignal_ROM_256x8 is
   subtype TDataWord is std_logic_vector(7 downto 0);
   type TROM is array (0 to 255) of TDataWord;
	-- Input Signal ROM
   constant c_memory: TROM := (
	"10000001",
	"10000101",
	"10001001",
	"10001110",
	"10010010",
	"10010110",
	"10011010",
	"10011111",
	"10100011",
	"10100111",
	"10101011",
	"10110000",
	"10110100",
	"10111000",
	"10111100",
	"11000000",
	"11000101",
	"11001001",
	"11001101",
	"11010001",
	"11010110",
	"11011010",
	"11011110",
	"11100010",
	"11100111",
	"11101011",
	"11101111",
	"11110011",
	"11111000",
	"11111100",
	"00000000",
	"00000100",
	"00001000",
	"00001101",
	"00010001",
	"00010101",
	"00011001",
	"00011110",
	"00100010",
	"00100110",
	"00101010",
	"00101111",
	"00110011",
	"00110111",
	"00111011",
	"01000000",
	"01000100",
	"01001000",
	"01001100",
	"01010000",
	"01010101",
	"01011001",
	"01011101",
	"01100001",
	"01100110",
	"01101010",
	"01101110",
	"01110010",
	"01110111",
	"01111011",
	"01111111",
	"01111011",
	"01110111",
	"01110010",
	"01101110",
	"01101010",
	"01100110",
	"01100001",
	"01011101",
	"01011001",
	"01010101",
	"01010000",
	"01001100",
	"01001000",
	"01000100",
	"01000000",
	"00111011",
	"00110111",
	"00110011",
	"00101111",
	"00101010",
	"00100110",
	"00100010",
	"00011110",
	"00011001",
	"00010101",
	"00010001",
	"00001101",
	"00001000",
	"00000100",
	"00000000",
	"11111100",
	"11111000",
	"11110011",
	"11101111",
	"11101011",
	"11100111",
	"11100010",
	"11011110",
	"11011010",
	"11010110",
	"11010001",
	"11001101",
	"11001001",
	"11000101",
	"11000000",
	"10111100",
	"10111000",
	"10110100",
	"10110000",
	"10101011",
	"10100111",
	"10100011",
	"10011111",
	"10011010",
	"10010110",
	"10010010",
	"10001110",
	"10001001",
	"10000101",
	"10000001",
	"10000101",
	"10001001",
	"10001110",
	"10010010",
	"10010110",
	"10011010",
	"10011111",
	"10100011",
	"10100111",
	"10101011",
	"10110000",
	"10110100",
	"10111000",
	"10111100",
	"11000000",
	"11000101",
	"11001001",
	"11001101",
	"11010001",
	"11010110",
	"11011010",
	"11011110",
	"11100010",
	"11100111",
	"11101011",
	"11101111",
	"11110011",
	"11111000",
	"11111100",
	"00000000",
	"00000100",
	"00001000",
	"00001101",
	"00010001",
	"00010101",
	"00011001",
	"00011110",
	"00100010",
	"00100110",
	"00101010",
	"00101111",
	"00110011",
	"00110111",
	"00111011",
	"00111111",
	"01000100",
	"01001000",
	"01001100",
	"01010000",
	"01010101",
	"01011001",
	"01011101",
	"01100001",
	"01100110",
	"01101010",
	"01101110",
	"01110010",
	"01110111",
	"01111011",
	"01111111",
	"01111011",
	"01110111",
	"01110010",
	"01101110",
	"01101010",
	"01100110",
	"01100001",
	"01011101",
	"01011001",
	"01010101",
	"01010000",
	"01001100",
	"01001000",
	"01000100",
	"01000000",
	"00111011",
	"00110111",
	"00110011",
	"00101111",
	"00101010",
	"00100110",
	"00100010",
	"00011110",
	"00011001",
	"00010101",
	"00010001",
	"00001101",
	"00001000",
	"00000100",
	"00000000",
	"11111100",
	"11111000",
	"11110011",
	"11101111",
	"11101011",
	"11100111",
	"11100010",
	"11011110",
	"11011010",
	"11010110",
	"11010001",
	"11001101",
	"11001001",
	"11000101",
	"11000001",
	"10111100",
	"10111000",
	"10110100",
	"10110000",
	"10101011",
	"10100111",
	"10100011",
	"10011111",
	"10011010",
	"10010110",
	"10010010",
	"10001110",
	"10001001",
	"10000101",
	"10000001",
	"10000101",
	"10001001",
	"10001110",
	"10010010",
	"10010110",
	"10011010",
	"10011111",
	"10100011",
	"10100111",
	"10101011",
	"10110000",
	"10110100",
	"10111000",
	"10111100",
	"11000000"
	);

begin
   dataOut <= c_memory(to_integer(unsigned(address)));
end Behavioral;
