-- Inclua as bibliotecas e os pacotes necessários
entity Adder4 is
 port(a, b  : in std_logic_vector(3 downto 0);
		cin 	: in std_logic;
		s 		: out std_logic_vector(3 downto 0);
		cout  : out std_logic);

end Adder4;

architecture Structural of Adder4 is

 -- Declare um sinal interno (carryOut) do tipo std_logic_vector (de
 -- C bits) que interligará os bits de carry dos somadores entre si
begin
	bit0: entity work.FullAdder(Behavioral)
			 port map(a => a(0),
						 b => b(0),
						 cin => cin,
						 s => s(0),
						 cout => carryOut(0));
-- complete para os restantes bits (1 a 3)
end Structural; 